library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity xor_gate is
port(a, b: in std_logic;
	  output: out std_logic);
end xor_gate;

architecture Behavioral of xor_gate is
begin

process (a, b)
begin
	if (a = b) then 
		output <= '0';
	else 
		output <= '1';
	end if;
end process;

end Behavioral;